package master_agent_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "master_seq_item.sv"
	`include "master_sequencer.sv"
	`include "master_sequence.sv"
	`include "master_agt_cfg.sv"
	`include "master_driver.sv"
	`include "master_monitor.sv"
	`include "master_agent.sv"
	`include "master_agt_top.sv"

endpackage: master_agent_pkg
