package slave_agent_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "slave_seq_item.sv"
	`include "slave_sequencer.sv"
	`include "slave_sequence.sv"
	`include "slave_agt_cfg.sv"
	`include "slave_driver.sv"
	`include "slave_monitor.sv"
	`include "slave_agent.sv"
	`include "slave_agt_top.sv"

endpackage: slave_agent_pkg
