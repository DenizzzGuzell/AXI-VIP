package axi_test_pkg;

	import uvm_pkg::*;
	import env_pkg::*;

	`include "uvm_macros.svh"
	`include "../master_agt_top/master_agt_cfg.sv"
	`include "../slave_agt_top/slave_agt_cfg.sv"
	`include "axi_test.sv"


endpackage
